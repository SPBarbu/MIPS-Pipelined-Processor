library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity processor is
end processor;

architecture behavior of processor is
begin

end;