library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity EX_stage is
end EX_stage;

architecture behavior of EX_stage is
begin

end;