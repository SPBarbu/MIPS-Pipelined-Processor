library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ID_stage is
end ID_stage;

architecture behavior of ID_stage is
begin

end;