library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IF_stage is
end IF_stage;

architecture behavior of IF_stage is
begin

end;