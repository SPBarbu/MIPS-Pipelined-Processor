library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WB_stage is
end WB_stage;

architecture behavior of WB_stage is
begin

end;