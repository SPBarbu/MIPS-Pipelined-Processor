library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MEM_stage is
end MEM_stage;

architecture behavior of MEM_stage is
begin

end;